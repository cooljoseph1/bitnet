module stoch_grad_tb();

    integer i;
    integer j;
    logic [12:0] k;
  logic rst_in = 0;
  logic clk_in = 0;

  localparam W_SIZE = 256;
  logic [W_SIZE-1:0] g_in = 0;
  logic [W_SIZE-1:0] g_out;

  stoch_grad #(
    .W_SIZE(W_SIZE)
  ) stoch_grad_test(
    .clk_in(clk_in),
    .rst_in(rst_in),
    .flip_weight_in(g_in),
    .flip_weight_out(g_out)
  );

  always begin
      #5;
      clk_in = !clk_in;
  end

  
  initial begin
    $dumpfile("stoch_grad.vcd"); //file to store value change dump (vcd)
    $dumpvars(1,stoch_grad_test);
    $display("\n--------\nStarting Simulation!");
    
    rst_in = 1;
    #10;
    rst_in = 0;
    #10;
    for (i=0; i<W_SIZE; i = i+1)begin
      k = 13'b1_1111_1111_1111;
      for(j=0; j < 8; j = j+1)begin
        k ^= 13'b1 << ((i * i * i * 17 + i * j * 19) % 13);
      end
      $display((k | 13'b1_0000_0000_0000));
    end

    #10
    
    g_in = 256'b110_100_1_100_1100_11_1101_1011_1010_1100_1010_1000_101_0_11_1101_1110_1001_110_1110_111_100_1110_1110_1011_1000_11_111_111_1110_101_110_100_1101_1110_1111_1111_110_101_1010_101_1111_101_110_1100_1001_1000_10_100_101_1000_1110_1_1110_11_101_1101_1000_100_1000_1101_1_1011_111_11_0_1101_1_110_11_0_1_11_1100_1001_1110_1001_11_1000_10_1010_1000_1101_1_1010_11_1_1_1000_10_110_10_1_1001_10_1011_100_1010_0_1001_1101_1010_11_1111_1011_1000_11_110_1110_1111_101_11_1001_11_1110_11_10_11_1_101_1101_1_1111_0_0_111_0_1_1101_100_1110_1001_1110_1_0_111_1101_110_100_1000_1000_11_111_1010_1_1000_1010_110_1_1111_1001_101_1_101_1101_1010_1000_1000_1110_1001_1010_1100_0_1001_111_1111_101_1_0_1110_1011_1111_1100_110_1111_111_1001_110_1010_100_100_1000_100_1101_1101_100_1011_1010_0_1111_111_0_110_1010_0_101_1010_10_111_1011_1000_110_1111_1010_1110_111_10_1111_1110_1001_1000_1100_1110_1100_1111_101_1_1111_10_10_1000_101_0_10_1110_1011_1000_1110_1101_1110_0_1011_1110_1110_11_1_1010_1010_0_111_1000_1010_1010_1_100_110_1001_0_1110_111_101_101_0_1000_1110_1011;
    $display(g_in);
    #10;
    #10;
    #10;
    #10;
    #10;
    $finish;
  end
endmodule // stoch_grad_tb