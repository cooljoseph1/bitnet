typedef enum bit [3:0] {RECV=0, SEND=1, READ=2, WRITE=3} op;